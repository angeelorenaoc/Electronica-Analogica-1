Rectificador

VP 1 0 SIN (0 170 60HZ  0 0 0)
L1 2 0 722.4M
L2 3 0 5M

KTRANS L1 L2 0.9999

D1 3 4 D1N4004
D2 5 0 D1N4004
D3 5 3 D1N4004
D4 0 4 D1N4004
RP 1 2 5U
RL 4 5 1000

.lib diode.lib
.PROBE
.TRAN 35u 35m 0 35u
.END


