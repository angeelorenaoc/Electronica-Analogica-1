Circuito de polarizaci�n de BJT
VCC 1 0 DC 12
RC 1 2 47K
R1 1 3 189.09447K
Q1 2 3 4 QNPN
RE 4 0 1.88071k
R2 3 0 20.8842182k
C1 5 3 10U
RSIG 5 7 50
V1 5 0 SIN(0 100m 5KHz 0 0 0)
C2 2 6 10U
RL 6 0 47K

.MODEL QNPN NPN (BF=100 VA=100)
.OP
.AC DEC 5000 1 10MEG
.PROBE
.END